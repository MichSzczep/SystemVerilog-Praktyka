// interface between DUT and TB


interface Counter_intface;
  logic CLK, reset, chnge;
  logic [3:0] load, out;
endinterface
